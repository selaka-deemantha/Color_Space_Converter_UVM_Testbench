package test_pkg;

    import uvm_pkg::*;  
    `include "uvm_macros.svh"

    import agent_pkg::*;
    import env_pkg::*;

    `include    "test.svh"

endpackage: test_pkg