package agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"



    `include "agent_config.svh"
    
    `include "seq_item.svh"
    `include "seq_item_in.svh"
    `include "seq_item_out.svh"
    `include "sequence_m.svh"

    `include "master_driver.svh"

    `include "master_monitor.svh"
    `include "slave_monitor.svh"

    `include "master_agent.svh"
    `include "slave_agent.svh"



endpackage: agent_pkg

