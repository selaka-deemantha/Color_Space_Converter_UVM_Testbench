package analysis_components_pkg;
    import      uvm_pkg::*;
    `include    "uvm_macros.svh"

    import      agent_pkg::*;

    `include    "checker_m.svh"
    `include    "predictor.svh"
    `include    "analysis_config.svh"
    
endpackage: analysis_components_pkg


