package env_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"


    import agent_pkg::*;
    import analysis_components_pkg::*;
    
    `include "env_config.svh"
    `include "env.svh"
    
endpackage: env_pkg